`timescale 1ns / 1ps

module rom_memory #(
    parameter SIZE_BYTES = 16384,
    parameter BASE_ADDR = 32'h80000000
)(
    input clk,
    input rst_n,
    
    input         mem_valid,
    output        mem_ready,
    input  [31:0] mem_addr,
    input  [31:0] mem_wdata,
    input  [3:0]  mem_wstrb,
    output [31:0] mem_rdata
);

    localparam SIZE_WORDS = SIZE_BYTES / 4;
    localparam ADDR_BITS = $clog2(SIZE_WORDS);

    // ROM storage
    reg [31:0] rom_data [0:SIZE_WORDS-1];

    // Address calculation
    wire [ADDR_BITS-1:0] word_addr = (mem_addr - BASE_ADDR) >> 2;
    
    // ROM is always ready for reads, ignores writes
    assign mem_ready = mem_valid;
    
    // Read data
    assign mem_rdata = mem_valid ? rom_data[word_addr] : 32'h0;

    // Initialize ROM with matrix test program
    integer i;
    initial begin
        // Initialize all locations to NOP (addi x0, x0, 0)
        for (i = 0; i < SIZE_WORDS; i = i + 1) begin
            rom_data[i] = 32'h00000013; // NOP instruction
        end
        
        // Load compiled program
        rom_data[   0] = 32'h00003117;  // 0x80000000
        rom_data[   1] = 32'h20010113;  // 0x80000004
        rom_data[   2] = 32'h132000ef;  // 0x80000008
        rom_data[   3] = 32'h00003297;  // 0x8000000c
        rom_data[   4] = 32'h1f428293;  // 0x80000010
        rom_data[   5] = 32'hb0234305;  // 0x80000014
        rom_data[   6] = 32'ha0010062;  // 0x80000018
        rom_data[   7] = 32'he4261101;  // 0x8000001c
        rom_data[   8] = 32'h8493e04a;  // 0x80000020
        rom_data[   9] = 32'h89130045;  // 0x80000024
        rom_data[  10] = 32'h85aa0145;  // 0x80000028
        rom_data[  11] = 32'h00001517;  // 0x8000002c
        rom_data[  12] = 32'hb0450513;  // 0x80000030
        rom_data[  13] = 32'he822ec06;  // 0x80000034
        rom_data[  14] = 32'h7cc000ef;  // 0x80000038
        rom_data[  15] = 32'h00001517;  // 0x8000003c
        rom_data[  16] = 32'hb0450513;  // 0x80000040
        rom_data[  17] = 32'h7c0000ef;  // 0x80000044
        rom_data[  18] = 32'hffc4c583;  // 0x80000048
        rom_data[  19] = 32'hffc48413;  // 0x8000004c
        rom_data[  20] = 32'h00001517;  // 0x80000050
        rom_data[  21] = 32'haf850513;  // 0x80000054
        rom_data[  22] = 32'h7ac000ef;  // 0x80000058
        rom_data[  23] = 32'h15170405;  // 0x8000005c
        rom_data[  24] = 32'h05130000;  // 0x80000060
        rom_data[  25] = 32'h0363afa5;  // 0x80000064
        rom_data[  26] = 32'h00ef0294;  // 0x80000068
        rom_data[  27] = 32'h458379a0;  // 0x8000006c
        rom_data[  28] = 32'h15170004;  // 0x80000070
        rom_data[  29] = 32'h05130000;  // 0x80000074
        rom_data[  30] = 32'h0405ad65;  // 0x80000078
        rom_data[  31] = 32'h788000ef;  // 0x8000007c
        rom_data[  32] = 32'h00001517;  // 0x80000080
        rom_data[  33] = 32'had850513;  // 0x80000084
        rom_data[  34] = 32'hfe9411e3;  // 0x80000088
        rom_data[  35] = 32'h00001517;  // 0x8000008c
        rom_data[  36] = 32'hac450513;  // 0x80000090
        rom_data[  37] = 32'h00440493;  // 0x80000094
        rom_data[  38] = 32'h24d000ef;  // 0x80000098
        rom_data[  39] = 32'hfb2490e3;  // 0x8000009c
        rom_data[  40] = 32'h644260e2;  // 0x800000a0
        rom_data[  41] = 32'h690264a2;  // 0x800000a4
        rom_data[  42] = 32'h80826105;  // 0x800000a8
        rom_data[  43] = 32'he4261101;  // 0x800000ac
        rom_data[  44] = 32'h8493e04a;  // 0x800000b0
        rom_data[  45] = 32'h89130105;  // 0x800000b4
        rom_data[  46] = 32'h85aa0505;  // 0x800000b8
        rom_data[  47] = 32'h00001517;  // 0x800000bc
        rom_data[  48] = 32'ha7450513;  // 0x800000c0
        rom_data[  49] = 32'he822ec06;  // 0x800000c4
        rom_data[  50] = 32'h73c000ef;  // 0x800000c8
        rom_data[  51] = 32'h00001517;  // 0x800000cc
        rom_data[  52] = 32'ha7450513;  // 0x800000d0
        rom_data[  53] = 32'h730000ef;  // 0x800000d4
        rom_data[  54] = 32'hff04a583;  // 0x800000d8
        rom_data[  55] = 32'hff048413;  // 0x800000dc
        rom_data[  56] = 32'h00001517;  // 0x800000e0
        rom_data[  57] = 32'ha8050513;  // 0x800000e4
        rom_data[  58] = 32'h71c000ef;  // 0x800000e8
        rom_data[  59] = 32'h15170411;  // 0x800000ec
        rom_data[  60] = 32'h05130000;  // 0x800000f0
        rom_data[  61] = 32'h0263a6a5;  // 0x800000f4
        rom_data[  62] = 32'h00ef0294;  // 0x800000f8
        rom_data[  63] = 32'h400c70a0;  // 0x800000fc
        rom_data[  64] = 32'h00001517;  // 0x80000100
        rom_data[  65] = 32'ha6050513;  // 0x80000104
        rom_data[  66] = 32'h00ef0411;  // 0x80000108
        rom_data[  67] = 32'h15176fa0;  // 0x8000010c
        rom_data[  68] = 32'h05130000;  // 0x80000110
        rom_data[  69] = 32'h12e3a4a5;  // 0x80000114
        rom_data[  70] = 32'h1517fe94;  // 0x80000118
        rom_data[  71] = 32'h05130000;  // 0x8000011c
        rom_data[  72] = 32'h0493a365;  // 0x80000120
        rom_data[  73] = 32'h00ef0104;  // 0x80000124
        rom_data[  74] = 32'h91e31bf0;  // 0x80000128
        rom_data[  75] = 32'h60e2fb24;  // 0x8000012c
        rom_data[  76] = 32'h64a26442;  // 0x80000130
        rom_data[  77] = 32'h61056902;  // 0x80000134
        rom_data[  78] = 32'h71718082;  // 0x80000138
        rom_data[  79] = 32'h00001517;  // 0x8000013c
        rom_data[  80] = 32'ha3c50513;  // 0x80000140
        rom_data[  81] = 32'he94af506;  // 0x80000144
        rom_data[  82] = 32'h19d000ef;  // 0x80000148
        rom_data[  83] = 32'h00001517;  // 0x8000014c
        rom_data[  84] = 32'ha5450513;  // 0x80000150
        rom_data[  85] = 32'h191000ef;  // 0x80000154
        rom_data[  86] = 32'h2ba000ef;  // 0x80000158
        rom_data[  87] = 32'h2a051063;  // 0x8000015c
        rom_data[  88] = 32'h84aaed26;  // 0x80000160
        rom_data[  89] = 32'h00001517;  // 0x80000164
        rom_data[  90] = 32'ha9450513;  // 0x80000168
        rom_data[  91] = 32'he54ef122;  // 0x8000016c
        rom_data[  92] = 32'hfcd6e152;  // 0x80000170
        rom_data[  93] = 32'h00eff8da;  // 0x80000174
        rom_data[  94] = 32'h059316f0;  // 0x80000178
        rom_data[  95] = 32'h051300f1;  // 0x8000017c
        rom_data[  96] = 32'h00ef00e1;  // 0x80000180
        rom_data[  97] = 32'hed0d5b80;  // 0x80000184
        rom_data[  98] = 32'h00e14783;  // 0x80000188
        rom_data[  99] = 32'h00001597;  // 0x8000018c
        rom_data[ 100] = 32'h9e458593;  // 0x80000190
        rom_data[ 101] = 32'h1597c789;  // 0x80000194
        rom_data[ 102] = 32'h85930000;  // 0x80000198
        rom_data[ 103] = 32'h47839d25;  // 0x8000019c
        rom_data[ 104] = 32'h161700f1;  // 0x800001a0
        rom_data[ 105] = 32'h06130000;  // 0x800001a4
        rom_data[ 106] = 32'hc7899ce6;  // 0x800001a8
        rom_data[ 107] = 32'h00001617;  // 0x800001ac
        rom_data[ 108] = 32'h9bc60613;  // 0x800001b0
        rom_data[ 109] = 32'h00001517;  // 0x800001b4
        rom_data[ 110] = 32'ha6c50513;  // 0x800001b8
        rom_data[ 111] = 32'h648000ef;  // 0x800001bc
        rom_data[ 112] = 32'h00001417;  // 0x800001c0
        rom_data[ 113] = 32'he8040413;  // 0x800001c4
        rom_data[ 114] = 32'h4a814901;  // 0x800001c8
        rom_data[ 115] = 32'h36034b41;  // 0x800001cc
        rom_data[ 116] = 32'h2485fd84;  // 0x800001d0
        rom_data[ 117] = 32'h151785a6;  // 0x800001d4
        rom_data[ 118] = 32'h05130000;  // 0x800001d8
        rom_data[ 119] = 32'h00efa725;  // 0x800001dc
        rom_data[ 120] = 32'h0a136260;  // 0x800001e0
        rom_data[ 121] = 32'h0993fe04;  // 0x800001e4
        rom_data[ 122] = 32'h6689ff04;  // 0x800001e8
        rom_data[ 123] = 32'h181085ce;  // 0x800001ec
        rom_data[ 124] = 32'h86938552;  // 0x800001f0
        rom_data[ 125] = 32'h00ef7106;  // 0x800001f4
        rom_data[ 126] = 32'h181041a0;  // 0x800001f8
        rom_data[ 127] = 32'h176385a2;  // 0x800001fc
        rom_data[ 128] = 32'h47811605;  // 0x80000200
        rom_data[ 129] = 32'h00f606b3;  // 0x80000204
        rom_data[ 130] = 32'h00f58733;  // 0x80000208
        rom_data[ 131] = 32'h43184294;  // 0x8000020c
        rom_data[ 132] = 32'h98630791;  // 0x80000210
        rom_data[ 133] = 32'h97e316e6;  // 0x80000214
        rom_data[ 134] = 32'h0641ff67;  // 0x80000218
        rom_data[ 135] = 32'h05c1189c;  // 0x8000021c
        rom_data[ 136] = 32'hfef611e3;  // 0x80000220
        rom_data[ 137] = 32'h151785a6;  // 0x80000224
        rom_data[ 138] = 32'h05130000;  // 0x80000228
        rom_data[ 139] = 32'h00efcba5;  // 0x8000022c
        rom_data[ 140] = 32'h2a855d60;  // 0x80000230
        rom_data[ 141] = 32'h00ef4529;  // 0x80000234
        rom_data[ 142] = 32'h478d0930;  // 0x80000238
        rom_data[ 143] = 32'h06840413;  // 0x8000023c
        rom_data[ 144] = 32'hf8f497e3;  // 0x80000240
        rom_data[ 145] = 32'h00001517;  // 0x80000244
        rom_data[ 146] = 32'ha5c50513;  // 0x80000248
        rom_data[ 147] = 32'h099000ef;  // 0x8000024c
        rom_data[ 148] = 32'h151785a6;  // 0x80000250
        rom_data[ 149] = 32'h05130000;  // 0x80000254
        rom_data[ 150] = 32'h00efa665;  // 0x80000258
        rom_data[ 151] = 32'h85d65aa0;  // 0x8000025c
        rom_data[ 152] = 32'h00001517;  // 0x80000260
        rom_data[ 153] = 32'ha7050513;  // 0x80000264
        rom_data[ 154] = 32'h59c000ef;  // 0x80000268
        rom_data[ 155] = 32'h151785ca;  // 0x8000026c
        rom_data[ 156] = 32'h05130000;  // 0x80000270
        rom_data[ 157] = 32'h00efa725;  // 0x80000274
        rom_data[ 158] = 32'hf7d358e0;  // 0x80000278
        rom_data[ 159] = 32'h1797d00a;  // 0x8000027c
        rom_data[ 160] = 32'ha6870000;  // 0x80000280
        rom_data[ 161] = 32'h1797f6a7;  // 0x80000284
        rom_data[ 162] = 32'ha7070000;  // 0x80000288
        rom_data[ 163] = 32'h1517f667;  // 0x8000028c
        rom_data[ 164] = 32'h05130000;  // 0x80000290
        rom_data[ 165] = 32'hf7d3a625;  // 0x80000294
        rom_data[ 166] = 32'hf7d318d7;  // 0x80000298
        rom_data[ 167] = 32'h87d310e7;  // 0x8000029c
        rom_data[ 168] = 32'h85d34207;  // 0x800002a0
        rom_data[ 169] = 32'h00efe207;  // 0x800002a4
        rom_data[ 170] = 32'h116355e0;  // 0x800002a8
        rom_data[ 171] = 32'h15171209;  // 0x800002ac
        rom_data[ 172] = 32'h05130000;  // 0x800002b0
        rom_data[ 173] = 32'h00efa5a5;  // 0x800002b4
        rom_data[ 174] = 32'h151702f0;  // 0x800002b8
        rom_data[ 175] = 32'h05130000;  // 0x800002bc
        rom_data[ 176] = 32'h00efa965;  // 0x800002c0
        rom_data[ 177] = 32'h17970230;  // 0x800002c4
        rom_data[ 178] = 32'h87930000;  // 0x800002c8
        rom_data[ 179] = 32'hb603d527;  // 0x800002cc
        rom_data[ 180] = 32'hb6831387;  // 0x800002d0
        rom_data[ 181] = 32'hb7031407;  // 0x800002d4
        rom_data[ 182] = 32'hb7831487;  // 0x800002d8
        rom_data[ 183] = 32'h15171507;  // 0x800002dc
        rom_data[ 184] = 32'h05130000;  // 0x800002e0
        rom_data[ 185] = 32'he832a9a5;  // 0x800002e4
        rom_data[ 186] = 32'hf03aec36;  // 0x800002e8
        rom_data[ 187] = 32'h00eff43e;  // 0x800002ec
        rom_data[ 188] = 32'h080c7f60;  // 0x800002f0
        rom_data[ 189] = 32'h00001517;  // 0x800002f4
        rom_data[ 190] = 32'hab450513;  // 0x800002f8
        rom_data[ 191] = 32'hd21ff0ef;  // 0x800002fc
        rom_data[ 192] = 32'h1517100c;  // 0x80000300
        rom_data[ 193] = 32'h05130000;  // 0x80000304
        rom_data[ 194] = 32'hf0efabe5;  // 0x80000308
        rom_data[ 195] = 32'h66b1d13f;  // 0x8000030c
        rom_data[ 196] = 32'h0808100c;  // 0x80000310
        rom_data[ 197] = 32'h86931810;  // 0x80000314
        rom_data[ 198] = 32'h00ef3506;  // 0x80000318
        rom_data[ 199] = 32'he5692f60;  // 0x8000031c
        rom_data[ 200] = 32'h00001517;  // 0x80000320
        rom_data[ 201] = 32'hab850513;  // 0x80000324
        rom_data[ 202] = 32'h7bc000ef;  // 0x80000328
        rom_data[ 203] = 32'h1517180c;  // 0x8000032c
        rom_data[ 204] = 32'h05130000;  // 0x80000330
        rom_data[ 205] = 32'hf0efada5;  // 0x80000334
        rom_data[ 206] = 32'h0593d77f;  // 0x80000338
        rom_data[ 207] = 32'h15173e80;  // 0x8000033c
        rom_data[ 208] = 32'h05130000;  // 0x80000340
        rom_data[ 209] = 32'h00efae25;  // 0x80000344
        rom_data[ 210] = 32'h15174be0;  // 0x80000348
        rom_data[ 211] = 32'h05130000;  // 0x8000034c
        rom_data[ 212] = 32'h00efaee5;  // 0x80000350
        rom_data[ 213] = 32'h740a7920;  // 0x80000354
        rom_data[ 214] = 32'h69aa64ea;  // 0x80000358
        rom_data[ 215] = 32'h7ae66a0a;  // 0x8000035c
        rom_data[ 216] = 32'h70aa7b46;  // 0x80000360
        rom_data[ 217] = 32'h694a854a;  // 0x80000364
        rom_data[ 218] = 32'h8082614d;  // 0x80000368
        rom_data[ 219] = 32'h3f4000ef;  // 0x8000036c
        rom_data[ 220] = 32'h151785aa;  // 0x80000370
        rom_data[ 221] = 32'h05130000;  // 0x80000374
        rom_data[ 222] = 32'h00ef8fe5;  // 0x80000378
        rom_data[ 223] = 32'h290548a0;  // 0x8000037c
        rom_data[ 224] = 32'h85a6bd6d;  // 0x80000380
        rom_data[ 225] = 32'h00001517;  // 0x80000384
        rom_data[ 226] = 32'hb7c50513;  // 0x80000388
        rom_data[ 227] = 32'h478000ef;  // 0x8000038c
        rom_data[ 228] = 32'h151785d2;  // 0x80000390
        rom_data[ 229] = 32'h05130000;  // 0x80000394
        rom_data[ 230] = 32'hf0efb8e5;  // 0x80000398
        rom_data[ 231] = 32'h85cec83f;  // 0x8000039c
        rom_data[ 232] = 32'h00001517;  // 0x800003a0
        rom_data[ 233] = 32'hb9050513;  // 0x800003a4
        rom_data[ 234] = 32'hc75ff0ef;  // 0x800003a8
        rom_data[ 235] = 32'h151785a2;  // 0x800003ac
        rom_data[ 236] = 32'h05130000;  // 0x800003b0
        rom_data[ 237] = 32'hf0efb925;  // 0x800003b4
        rom_data[ 238] = 32'h180ccf7f;  // 0x800003b8
        rom_data[ 239] = 32'h00001517;  // 0x800003bc
        rom_data[ 240] = 32'hb9450513;  // 0x800003c0
        rom_data[ 241] = 32'hce9ff0ef;  // 0x800003c4
        rom_data[ 242] = 32'hb5ad2905;  // 0x800003c8
        rom_data[ 243] = 32'h00001517;  // 0x800003cc
        rom_data[ 244] = 32'hacc50513;  // 0x800003d0
        rom_data[ 245] = 32'h710000ef;  // 0x800003d4
        rom_data[ 246] = 32'h740a597d;  // 0x800003d8
        rom_data[ 247] = 32'h69aa64ea;  // 0x800003dc
        rom_data[ 248] = 32'h7ae66a0a;  // 0x800003e0
        rom_data[ 249] = 32'hbfb57b46;  // 0x800003e4
        rom_data[ 250] = 32'h378000ef;  // 0x800003e8
        rom_data[ 251] = 32'h151785aa;  // 0x800003ec
        rom_data[ 252] = 32'h05130000;  // 0x800003f0
        rom_data[ 253] = 32'h00efa8a5;  // 0x800003f4
        rom_data[ 254] = 32'hbfb140e0;  // 0x800003f8
        rom_data[ 255] = 32'h364000ef;  // 0x800003fc
        rom_data[ 256] = 32'h051785aa;  // 0x80000400
        rom_data[ 257] = 32'h05130000;  // 0x80000404
        rom_data[ 258] = 32'h00ef7c65;  // 0x80000408
        rom_data[ 259] = 32'h597d3fa0;  // 0x8000040c
        rom_data[ 260] = 32'h07b7bf89;  // 0x80000410
        rom_data[ 261] = 32'h47091000;  // 0x80000414
        rom_data[ 262] = 32'hc3981141;  // 0x80000418
        rom_data[ 263] = 32'h47b2c602;  // 0x8000041c
        rom_data[ 264] = 32'h06300713;  // 0x80000420
        rom_data[ 265] = 32'h00f76963;  // 0x80000424
        rom_data[ 266] = 32'h47b20001;  // 0x80000428
        rom_data[ 267] = 32'hc63e2785;  // 0x8000042c
        rom_data[ 268] = 32'h7be347b2;  // 0x80000430
        rom_data[ 269] = 32'h07b7fef7;  // 0x80000434
        rom_data[ 270] = 32'ha0231000;  // 0x80000438
        rom_data[ 271] = 32'hc4020007;  // 0x8000043c
        rom_data[ 272] = 32'h071347a2;  // 0x80000440
        rom_data[ 273] = 32'h69630630;  // 0x80000444
        rom_data[ 274] = 32'h000100f7;  // 0x80000448
        rom_data[ 275] = 32'h278547a2;  // 0x8000044c
        rom_data[ 276] = 32'h47a2c43e;  // 0x80000450
        rom_data[ 277] = 32'hfef77be3;  // 0x80000454
        rom_data[ 278] = 32'h000407b7;  // 0x80000458
        rom_data[ 279] = 32'h10000737;  // 0x8000045c
        rom_data[ 280] = 32'h40478793;  // 0x80000460
        rom_data[ 281] = 32'h0721c71c;  // 0x80000464
        rom_data[ 282] = 32'h15634318;  // 0x80000468
        rom_data[ 283] = 32'h450100f7;  // 0x8000046c
        rom_data[ 284] = 32'h80820141;  // 0x80000470
        rom_data[ 285] = 32'hbfed5575;  // 0x80000474
        rom_data[ 286] = 32'h100007b7;  // 0x80000478
        rom_data[ 287] = 32'h810543c8;  // 0x8000047c
        rom_data[ 288] = 32'h45138905;  // 0x80000480
        rom_data[ 289] = 32'h80820015;  // 0x80000484
        rom_data[ 290] = 32'h100007b7;  // 0x80000488
        rom_data[ 291] = 32'h890543c8;  // 0x8000048c
        rom_data[ 292] = 32'h07b78082;  // 0x80000490
        rom_data[ 293] = 32'h07911000;  // 0x80000494
        rom_data[ 294] = 32'h8b89439c;  // 0x80000498
        rom_data[ 295] = 32'h0637eb9d;  // 0x8000049c
        rom_data[ 296] = 32'h05111000;  // 0x800004a0
        rom_data[ 297] = 32'h10060613;  // 0x800004a4
        rom_data[ 298] = 32'h48414581;  // 0x800004a8
        rom_data[ 299] = 32'hffc50793;  // 0x800004ac
        rom_data[ 300] = 32'hc6838732;  // 0x800004b0
        rom_data[ 301] = 32'h07850007;  // 0x800004b4
        rom_data[ 302] = 32'h2e230711;  // 0x800004b8
        rom_data[ 303] = 32'h9ae3fed7;  // 0x800004bc
        rom_data[ 304] = 32'h2591fea7;  // 0x800004c0
        rom_data[ 305] = 32'h85130641;  // 0x800004c4
        rom_data[ 306] = 32'h91e30047;  // 0x800004c8
        rom_data[ 307] = 32'h4501ff05;  // 0x800004cc
        rom_data[ 308] = 32'h55798082;  // 0x800004d0
        rom_data[ 309] = 32'h07b78082;  // 0x800004d4
        rom_data[ 310] = 32'h07911000;  // 0x800004d8
        rom_data[ 311] = 32'h8b89439c;  // 0x800004dc
        rom_data[ 312] = 32'h0637eb9d;  // 0x800004e0
        rom_data[ 313] = 32'h05111000;  // 0x800004e4
        rom_data[ 314] = 32'h20060613;  // 0x800004e8
        rom_data[ 315] = 32'h48414581;  // 0x800004ec
        rom_data[ 316] = 32'hffc50793;  // 0x800004f0
        rom_data[ 317] = 32'hc6838732;  // 0x800004f4
        rom_data[ 318] = 32'h07850007;  // 0x800004f8
        rom_data[ 319] = 32'h2e230711;  // 0x800004fc
        rom_data[ 320] = 32'h9ae3fed7;  // 0x80000500
        rom_data[ 321] = 32'h2591fea7;  // 0x80000504
        rom_data[ 322] = 32'h85130641;  // 0x80000508
        rom_data[ 323] = 32'h91e30047;  // 0x8000050c
        rom_data[ 324] = 32'h4501ff05;  // 0x80000510
        rom_data[ 325] = 32'h55798082;  // 0x80000514
        rom_data[ 326] = 32'h11418082;  // 0x80000518
        rom_data[ 327] = 32'he406e022;  // 0x8000051c
        rom_data[ 328] = 32'hf0ef842e;  // 0x80000520
        rom_data[ 329] = 32'he909f71f;  // 0x80000524
        rom_data[ 330] = 32'hf0ef8522;  // 0x80000528
        rom_data[ 331] = 32'he509fadf;  // 0x8000052c
        rom_data[ 332] = 32'h640260a2;  // 0x80000530
        rom_data[ 333] = 32'h80820141;  // 0x80000534
        rom_data[ 334] = 32'hbfdd5579;  // 0x80000538
        rom_data[ 335] = 32'h100007b7;  // 0x8000053c
        rom_data[ 336] = 32'h439c0791;  // 0x80000540
        rom_data[ 337] = 32'heb8d8b89;  // 0x80000544
        rom_data[ 338] = 32'h10000737;  // 0x80000548
        rom_data[ 339] = 32'h11414785;  // 0x8000054c
        rom_data[ 340] = 32'hc602c31c;  // 0x80000550
        rom_data[ 341] = 32'h474d47b2;  // 0x80000554
        rom_data[ 342] = 32'h00f76963;  // 0x80000558
        rom_data[ 343] = 32'h47b20001;  // 0x8000055c
        rom_data[ 344] = 32'hc63e2785;  // 0x80000560
        rom_data[ 345] = 32'h7be347b2;  // 0x80000564
        rom_data[ 346] = 32'h07b7fef7;  // 0x80000568
        rom_data[ 347] = 32'ha0231000;  // 0x8000056c
        rom_data[ 348] = 32'h45010007;  // 0x80000570
        rom_data[ 349] = 32'h80820141;  // 0x80000574
        rom_data[ 350] = 32'h80825579;  // 0x80000578
        rom_data[ 351] = 32'h10000637;  // 0x8000057c
        rom_data[ 352] = 32'h0611425c;  // 0x80000580
        rom_data[ 353] = 32'hef8d8b85;  // 0x80000584
        rom_data[ 354] = 32'h059b1141;  // 0x80000588
        rom_data[ 355] = 32'h4681fff5;  // 0x8000058c
        rom_data[ 356] = 32'hc6024725;  // 0x80000590
        rom_data[ 357] = 32'h696347b2;  // 0x80000594
        rom_data[ 358] = 32'h000100f7;  // 0x80000598
        rom_data[ 359] = 32'h278547b2;  // 0x8000059c
        rom_data[ 360] = 32'h47b2c63e;  // 0x800005a0
        rom_data[ 361] = 32'hfef77be3;  // 0x800005a4
        rom_data[ 362] = 32'h8b85421c;  // 0x800005a8
        rom_data[ 363] = 32'h2685e799;  // 0x800005ac
        rom_data[ 364] = 32'hfed5f1e3;  // 0x800005b0
        rom_data[ 365] = 32'h0141557d;  // 0x800005b4
        rom_data[ 366] = 32'h45018082;  // 0x800005b8
        rom_data[ 367] = 32'h80820141;  // 0x800005bc
        rom_data[ 368] = 32'h80824501;  // 0x800005c0
        rom_data[ 369] = 32'h100007b7;  // 0x800005c4
        rom_data[ 370] = 32'h439c0791;  // 0x800005c8
        rom_data[ 371] = 32'hcf9d8b85;  // 0x800005cc
        rom_data[ 372] = 32'h100008b7;  // 0x800005d0
        rom_data[ 373] = 32'h01050613;  // 0x800005d4
        rom_data[ 374] = 32'h30088893;  // 0x800005d8
        rom_data[ 375] = 32'h45814801;  // 0x800005dc
        rom_data[ 376] = 32'h06b34341;  // 0x800005e0
        rom_data[ 377] = 32'h8e890118;  // 0x800005e4
        rom_data[ 378] = 32'h873387aa;  // 0x800005e8
        rom_data[ 379] = 32'h431800f6;  // 0x800005ec
        rom_data[ 380] = 32'hae230791;  // 0x800005f0
        rom_data[ 381] = 32'h9ae3fee7;  // 0x800005f4
        rom_data[ 382] = 32'h2591fec7;  // 0x800005f8
        rom_data[ 383] = 32'h08410541;  // 0x800005fc
        rom_data[ 384] = 32'h01078613;  // 0x80000600
        rom_data[ 385] = 32'hfc659fe3;  // 0x80000604
        rom_data[ 386] = 32'h80824501;  // 0x80000608
        rom_data[ 387] = 32'h80825579;  // 0x8000060c
        rom_data[ 388] = 32'hf8227139;  // 0x80000610
        rom_data[ 389] = 32'hfc06f426;  // 0x80000614
        rom_data[ 390] = 32'h84b2e42e;  // 0x80000618
        rom_data[ 391] = 32'hf0ef8436;  // 0x8000061c
        rom_data[ 392] = 32'he561e75f;  // 0x80000620
        rom_data[ 393] = 32'hf0ef6522;  // 0x80000624
        rom_data[ 394] = 32'he161eb1f;  // 0x80000628
        rom_data[ 395] = 32'h100007b7;  // 0x8000062c
        rom_data[ 396] = 32'h07b743d4;  // 0x80000630
        rom_data[ 397] = 32'h8a891000;  // 0x80000634
        rom_data[ 398] = 32'h4705eacd;  // 0x80000638
        rom_data[ 399] = 32'hcc02c398;  // 0x8000063c
        rom_data[ 400] = 32'h474d47e2;  // 0x80000640
        rom_data[ 401] = 32'h00f76963;  // 0x80000644
        rom_data[ 402] = 32'h47e20001;  // 0x80000648
        rom_data[ 403] = 32'hcc3e2785;  // 0x8000064c
        rom_data[ 404] = 32'h7be347e2;  // 0x80000650
        rom_data[ 405] = 32'h07b7fef7;  // 0x80000654
        rom_data[ 406] = 32'ha0231000;  // 0x80000658
        rom_data[ 407] = 32'h86130007;  // 0x8000065c
        rom_data[ 408] = 32'h421c0047;  // 0x80000660
        rom_data[ 409] = 32'hfff4059b;  // 0x80000664
        rom_data[ 410] = 32'h8b854725;  // 0x80000668
        rom_data[ 411] = 32'hce02eb85;  // 0x8000066c
        rom_data[ 412] = 32'h696347f2;  // 0x80000670
        rom_data[ 413] = 32'h000100f7;  // 0x80000674
        rom_data[ 414] = 32'h278547f2;  // 0x80000678
        rom_data[ 415] = 32'h47f2ce3e;  // 0x8000067c
        rom_data[ 416] = 32'hfef77be3;  // 0x80000680
        rom_data[ 417] = 32'h8b85421c;  // 0x80000684
        rom_data[ 418] = 32'h2685eb91;  // 0x80000688
        rom_data[ 419] = 32'hfed5f1e3;  // 0x8000068c
        rom_data[ 420] = 32'h70e2557d;  // 0x80000690
        rom_data[ 421] = 32'h74a27442;  // 0x80000694
        rom_data[ 422] = 32'h80826121;  // 0x80000698
        rom_data[ 423] = 32'h100007b7;  // 0x8000069c
        rom_data[ 424] = 32'h439c0791;  // 0x800006a0
        rom_data[ 425] = 32'hc3b18b85;  // 0x800006a4
        rom_data[ 426] = 32'h10000337;  // 0x800006a8
        rom_data[ 427] = 32'h85938626;  // 0x800006ac
        rom_data[ 428] = 32'h03130104;  // 0x800006b0
        rom_data[ 429] = 32'h48813003;  // 0x800006b4
        rom_data[ 430] = 32'h4e414801;  // 0x800006b8
        rom_data[ 431] = 32'h006806b3;  // 0x800006bc
        rom_data[ 432] = 32'h87b28e91;  // 0x800006c0
        rom_data[ 433] = 32'h00f68733;  // 0x800006c4
        rom_data[ 434] = 32'h07914318;  // 0x800006c8
        rom_data[ 435] = 32'hfee7ae23;  // 0x800006cc
        rom_data[ 436] = 32'hfeb79ae3;  // 0x800006d0
        rom_data[ 437] = 32'h06412891;  // 0x800006d4
        rom_data[ 438] = 32'h05c10841;  // 0x800006d8
        rom_data[ 439] = 32'hffc890e3;  // 0x800006dc
        rom_data[ 440] = 32'h744270e2;  // 0x800006e0
        rom_data[ 441] = 32'h612174a2;  // 0x800006e4
        rom_data[ 442] = 32'h55798082;  // 0x800006e8
        rom_data[ 443] = 32'h07b7b75d;  // 0x800006ec
        rom_data[ 444] = 32'h47091000;  // 0x800006f0
        rom_data[ 445] = 32'hc3981141;  // 0x800006f4
        rom_data[ 446] = 32'h47b2c602;  // 0x800006f8
        rom_data[ 447] = 32'h06300713;  // 0x800006fc
        rom_data[ 448] = 32'h00f76963;  // 0x80000700
        rom_data[ 449] = 32'h47b20001;  // 0x80000704
        rom_data[ 450] = 32'hc63e2785;  // 0x80000708
        rom_data[ 451] = 32'h7be347b2;  // 0x8000070c
        rom_data[ 452] = 32'h07b7fef7;  // 0x80000710
        rom_data[ 453] = 32'ha0231000;  // 0x80000714
        rom_data[ 454] = 32'hc4020007;  // 0x80000718
        rom_data[ 455] = 32'h071347a2;  // 0x8000071c
        rom_data[ 456] = 32'h69630630;  // 0x80000720
        rom_data[ 457] = 32'h000100f7;  // 0x80000724
        rom_data[ 458] = 32'h278547a2;  // 0x80000728
        rom_data[ 459] = 32'h47a2c43e;  // 0x8000072c
        rom_data[ 460] = 32'hfef77be3;  // 0x80000730
        rom_data[ 461] = 32'h01414501;  // 0x80000734
        rom_data[ 462] = 32'h86aa8082;  // 0x80000738
        rom_data[ 463] = 32'hcd99c105;  // 0x8000073c
        rom_data[ 464] = 32'h100007b7;  // 0x80000740
        rom_data[ 465] = 32'h439c0791;  // 0x80000744
        rom_data[ 466] = 32'hd7134501;  // 0x80000748
        rom_data[ 467] = 32'h8b050017;  // 0x8000074c
        rom_data[ 468] = 32'h00e68023;  // 0x80000750
        rom_data[ 469] = 32'h80238b85;  // 0x80000754
        rom_data[ 470] = 32'h808200f5;  // 0x80000758
        rom_data[ 471] = 32'h80825575;  // 0x8000075c
        rom_data[ 472] = 32'h478d250d;  // 0x80000760
        rom_data[ 473] = 32'h00a7ed63;  // 0x80000764
        rom_data[ 474] = 32'h02051793;  // 0x80000768
        rom_data[ 475] = 32'h01d7d513;  // 0x8000076c
        rom_data[ 476] = 32'h00001797;  // 0x80000770
        rom_data[ 477] = 32'ha0078793;  // 0x80000774
        rom_data[ 478] = 32'h638897aa;  // 0x80000778
        rom_data[ 479] = 32'h15178082;  // 0x8000077c
        rom_data[ 480] = 32'h05130000;  // 0x80000780
        rom_data[ 481] = 32'h80828225;  // 0x80000784
        rom_data[ 482] = 32'h00001797;  // 0x80000788
        rom_data[ 483] = 32'h87878793;  // 0x8000078c
        rom_data[ 484] = 32'h0007b803;  // 0x80000790
        rom_data[ 485] = 32'h17976794;  // 0x80000794
        rom_data[ 486] = 32'hc7830000;  // 0x80000798
        rom_data[ 487] = 32'h713987a7;  // 0x8000079c
        rom_data[ 488] = 32'he836e442;  // 0x800007a0
        rom_data[ 489] = 32'h00f10c23;  // 0x800007a4
        rom_data[ 490] = 32'h1014c929;  // 0x800007a8
        rom_data[ 491] = 32'h8836872a;  // 0x800007ac
        rom_data[ 492] = 32'h77bb4501;  // 0x800007b0
        rom_data[ 493] = 32'h88ba02c7;  // 0x800007b4
        rom_data[ 494] = 32'h0805832a;  // 0x800007b8
        rom_data[ 495] = 32'h17822505;  // 0x800007bc
        rom_data[ 496] = 32'h978a9381;  // 0x800007c0
        rom_data[ 497] = 32'h0087c783;  // 0x800007c4
        rom_data[ 498] = 32'h02c7573b;  // 0x800007c8
        rom_data[ 499] = 32'hfef80fa3;  // 0x800007cc
        rom_data[ 500] = 32'hfec8f1e3;  // 0x800007d0
        rom_data[ 501] = 32'h00158613;  // 0x800007d4
        rom_data[ 502] = 32'h00d30733;  // 0x800007d8
        rom_data[ 503] = 32'h87ae961a;  // 0x800007dc
        rom_data[ 504] = 32'h00074683;  // 0x800007e0
        rom_data[ 505] = 32'h177d0785;  // 0x800007e4
        rom_data[ 506] = 32'hfed78fa3;  // 0x800007e8
        rom_data[ 507] = 32'hfec79ae3;  // 0x800007ec
        rom_data[ 508] = 32'h802395aa;  // 0x800007f0
        rom_data[ 509] = 32'h61210005;  // 0x800007f4
        rom_data[ 510] = 32'h80238082;  // 0x800007f8
        rom_data[ 511] = 32'h45010005;  // 0x800007fc
        rom_data[ 512] = 32'h80826121;  // 0x80000800
        rom_data[ 513] = 32'he5267115;  // 0x80000804
        rom_data[ 514] = 32'hed06e5be;  // 0x80000808
        rom_data[ 515] = 32'hf52efcce;  // 0x8000080c
        rom_data[ 516] = 32'hfd36f932;  // 0x80000810
        rom_data[ 517] = 32'he9c2e1ba;  // 0x80000814
        rom_data[ 518] = 32'h84aaedc6;  // 0x80000818
        rom_data[ 519] = 32'h00054503;  // 0x8000081c
        rom_data[ 520] = 32'he43e113c;  // 0x80000820
        rom_data[ 521] = 32'h1e050d63;  // 0x80000824
        rom_data[ 522] = 32'hf4d6f8d2;  // 0x80000828
        rom_data[ 523] = 32'hecdef0da;  // 0x8000082c
        rom_data[ 524] = 32'he922e8e2;  // 0x80000830
        rom_data[ 525] = 32'he4e6e14a;  // 0x80000834
        rom_data[ 526] = 32'h4981e0ea;  // 0x80000838
        rom_data[ 527] = 32'h02500a13;  // 0x8000083c
        rom_data[ 528] = 32'h07800a93;  // 0x80000840
        rom_data[ 529] = 32'h06200b13;  // 0x80000844
        rom_data[ 530] = 32'h1b974c55;  // 0x80000848
        rom_data[ 531] = 32'h8b930000;  // 0x8000084c
        rom_data[ 532] = 32'h8913946b;  // 0x80000850
        rom_data[ 533] = 32'h13630014;  // 0x80000854
        rom_data[ 534] = 32'hc7831745;  // 0x80000858
        rom_data[ 535] = 32'hef630014;  // 0x8000085c
        rom_data[ 536] = 32'h7a6300fa;  // 0x80000860
        rom_data[ 537] = 32'h879b12fb;  // 0x80000864
        rom_data[ 538] = 32'hf793f9d7;  // 0x80000868
        rom_data[ 539] = 32'h67630ff7;  // 0x8000086c
        rom_data[ 540] = 32'h078a00fc;  // 0x80000870
        rom_data[ 541] = 32'h439c97de;  // 0x80000874
        rom_data[ 542] = 32'h878297de;  // 0x80000878
        rom_data[ 543] = 32'h02500513;  // 0x8000087c
        rom_data[ 544] = 32'h248000ef;  // 0x80000880
        rom_data[ 545] = 32'h0014c503;  // 0x80000884
        rom_data[ 546] = 32'h00ef2989;  // 0x80000888
        rom_data[ 547] = 32'hc50323e0;  // 0x8000088c
        rom_data[ 548] = 32'h04930024;  // 0x80000890
        rom_data[ 549] = 32'hfd550019;  // 0x80000894
        rom_data[ 550] = 32'h60ea644a;  // 0x80000898
        rom_data[ 551] = 32'h7a46690a;  // 0x8000089c
        rom_data[ 552] = 32'h7b067aa6;  // 0x800008a0
        rom_data[ 553] = 32'h6c466be6;  // 0x800008a4
        rom_data[ 554] = 32'h6d066ca6;  // 0x800008a8
        rom_data[ 555] = 32'h854e64aa;  // 0x800008ac
        rom_data[ 556] = 32'h612d79e6;  // 0x800008b0
        rom_data[ 557] = 32'h67a28082;  // 0x800008b4
        rom_data[ 558] = 32'h07a14388;  // 0x800008b8
        rom_data[ 559] = 32'h0363e43e;  // 0x800008bc
        rom_data[ 560] = 32'h08001205;  // 0x800008c0
        rom_data[ 561] = 32'h464185a2;  // 0x800008c4
        rom_data[ 562] = 32'hec1ff0ef;  // 0x800008c8
        rom_data[ 563] = 32'hd1618d2a;  // 0x800008cc
        rom_data[ 564] = 32'h008d0cb3;  // 0x800008d0
        rom_data[ 565] = 32'h00044503;  // 0x800008d4
        rom_data[ 566] = 32'h00ef0405;  // 0x800008d8
        rom_data[ 567] = 32'h9be31ee0;  // 0x800008dc
        rom_data[ 568] = 32'hc503fe8c;  // 0x800008e0
        rom_data[ 569] = 32'h89bb0024;  // 0x800008e4
        rom_data[ 570] = 32'hb76501a9;  // 0x800008e8
        rom_data[ 571] = 32'h438867a2;  // 0x800008ec
        rom_data[ 572] = 32'he43e07a1;  // 0x800008f0
        rom_data[ 573] = 32'h0e050163;  // 0x800008f4
        rom_data[ 574] = 32'h85a20800;  // 0x800008f8
        rom_data[ 575] = 32'hf0ef4629;  // 0x800008fc
        rom_data[ 576] = 32'h8d2ae8bf;  // 0x80000900
        rom_data[ 577] = 32'h0cb3d549;  // 0x80000904
        rom_data[ 578] = 32'h4503008d;  // 0x80000908
        rom_data[ 579] = 32'h04050004;  // 0x8000090c
        rom_data[ 580] = 32'h1b8000ef;  // 0x80000910
        rom_data[ 581] = 32'hfe8c9be3;  // 0x80000914
        rom_data[ 582] = 32'h0024c503;  // 0x80000918
        rom_data[ 583] = 32'h01a989bb;  // 0x8000091c
        rom_data[ 584] = 32'h67a2bf8d;  // 0x80000920
        rom_data[ 585] = 32'h0007bc83;  // 0x80000924
        rom_data[ 586] = 32'he43e07a1;  // 0x80000928
        rom_data[ 587] = 32'h000cc503;  // 0x8000092c
        rom_data[ 588] = 32'hdd318466;  // 0x80000930
        rom_data[ 589] = 32'h194000ef;  // 0x80000934
        rom_data[ 590] = 32'h00144503;  // 0x80000938
        rom_data[ 591] = 32'hf97d0405;  // 0x8000093c
        rom_data[ 592] = 32'h4194043b;  // 0x80000940
        rom_data[ 593] = 32'h0024c503;  // 0x80000944
        rom_data[ 594] = 32'h013409bb;  // 0x80000948
        rom_data[ 595] = 32'h67a2b799;  // 0x8000094c
        rom_data[ 596] = 32'h07a14388;  // 0x80000950
        rom_data[ 597] = 32'h4e63e43e;  // 0x80000954
        rom_data[ 598] = 32'hc95d0805;  // 0x80000958
        rom_data[ 599] = 32'h85a20800;  // 0x8000095c
        rom_data[ 600] = 32'hf0ef4629;  // 0x80000960
        rom_data[ 601] = 32'h8d2ae27f;  // 0x80000964
        rom_data[ 602] = 32'h0cb3d11d;  // 0x80000968
        rom_data[ 603] = 32'h4503008d;  // 0x8000096c
        rom_data[ 604] = 32'h04050004;  // 0x80000970
        rom_data[ 605] = 32'h154000ef;  // 0x80000974
        rom_data[ 606] = 32'hfe8c9be3;  // 0x80000978
        rom_data[ 607] = 32'h0024c503;  // 0x8000097c
        rom_data[ 608] = 32'h01a989bb;  // 0x80000980
        rom_data[ 609] = 32'h67a2b739;  // 0x80000984
        rom_data[ 610] = 32'h43882985;  // 0x80000988
        rom_data[ 611] = 32'he43e07a1;  // 0x8000098c
        rom_data[ 612] = 32'h138000ef;  // 0x80000990
        rom_data[ 613] = 32'h8a63bded;  // 0x80000994
        rom_data[ 614] = 32'h071302a7;  // 0x80000998
        rom_data[ 615] = 32'h9fe302e0;  // 0x8000099c
        rom_data[ 616] = 32'hc503ece7;  // 0x800009a0
        rom_data[ 617] = 32'h07930024;  // 0x800009a4
        rom_data[ 618] = 32'h14e30310;  // 0x800009a8
        rom_data[ 619] = 32'hc703eef5;  // 0x800009ac
        rom_data[ 620] = 32'h07930034;  // 0x800009b0
        rom_data[ 621] = 32'h0b630660;  // 0x800009b4
        rom_data[ 622] = 32'h048906f7;  // 0x800009b8
        rom_data[ 623] = 32'h10c000ef;  // 0x800009bc
        rom_data[ 624] = 32'h0014c503;  // 0x800009c0
        rom_data[ 625] = 32'h89262985;  // 0x800009c4
        rom_data[ 626] = 32'h00efb5e9;  // 0x800009c8
        rom_data[ 627] = 32'hc5030fe0;  // 0x800009cc
        rom_data[ 628] = 32'h29850024;  // 0x800009d0
        rom_data[ 629] = 32'h0793bd7d;  // 0x800009d4
        rom_data[ 630] = 32'h18230300;  // 0x800009d8
        rom_data[ 631] = 32'h4d0500f1;  // 0x800009dc
        rom_data[ 632] = 32'hb7150800;  // 0x800009e0
        rom_data[ 633] = 32'h03000793;  // 0x800009e4
        rom_data[ 634] = 32'h00f11823;  // 0x800009e8
        rom_data[ 635] = 32'h08004d05;  // 0x800009ec
        rom_data[ 636] = 32'h0793b5c5;  // 0x800009f0
        rom_data[ 637] = 32'h053b02d0;  // 0x800009f4
        rom_data[ 638] = 32'h462940a0;  // 0x800009f8
        rom_data[ 639] = 32'h01110593;  // 0x800009fc
        rom_data[ 640] = 32'h00f10823;  // 0x80000a00
        rom_data[ 641] = 32'hd85ff0ef;  // 0x80000a04
        rom_data[ 642] = 32'h00150d1b;  // 0x80000a08
        rom_data[ 643] = 32'hbfb10800;  // 0x80000a0c
        rom_data[ 644] = 32'h03000793;  // 0x80000a10
        rom_data[ 645] = 32'h00f11823;  // 0x80000a14
        rom_data[ 646] = 32'h08004d05;  // 0x80000a18
        rom_data[ 647] = 32'h60eab7b9;  // 0x80000a1c
        rom_data[ 648] = 32'h64aa4981;  // 0x80000a20
        rom_data[ 649] = 32'h79e6854e;  // 0x80000a24
        rom_data[ 650] = 32'h8082612d;  // 0x80000a28
        rom_data[ 651] = 32'h071767a2;  // 0x80000a2c
        rom_data[ 652] = 32'h37070000;  // 0x80000a30
        rom_data[ 653] = 32'hfc6e7c27;  // 0x80000a34
        rom_data[ 654] = 32'h07a1239c;  // 0x80000a38
        rom_data[ 655] = 32'h9553e43e;  // 0x80000a3c
        rom_data[ 656] = 32'h8913c207;  // 0x80000a40
        rom_data[ 657] = 32'h06d30034;  // 0x80000a44
        rom_data[ 658] = 32'hf7d3d205;  // 0x80000a48
        rom_data[ 659] = 32'hf7d30ad7;  // 0x80000a4c
        rom_data[ 660] = 32'h97d312e7;  // 0x80000a50
        rom_data[ 661] = 32'h8dbec207;  // 0x80000a54
        rom_data[ 662] = 32'h04054963;  // 0x80000a58
        rom_data[ 663] = 32'h0800c121;  // 0x80000a5c
        rom_data[ 664] = 32'h462985a2;  // 0x80000a60
        rom_data[ 665] = 32'hd25ff0ef;  // 0x80000a64
        rom_data[ 666] = 32'hcd018d2a;  // 0x80000a68
        rom_data[ 667] = 32'h008d0cb3;  // 0x80000a6c
        rom_data[ 668] = 32'h00044503;  // 0x80000a70
        rom_data[ 669] = 32'h00ef0405;  // 0x80000a74
        rom_data[ 670] = 32'h9be30520;  // 0x80000a78
        rom_data[ 671] = 32'h89bbfe8c;  // 0x80000a7c
        rom_data[ 672] = 32'h051301a9;  // 0x80000a80
        rom_data[ 673] = 32'h00ef02e0;  // 0x80000a84
        rom_data[ 674] = 32'h851b0420;  // 0x80000a88
        rom_data[ 675] = 32'h00ef030d;  // 0x80000a8c
        rom_data[ 676] = 32'hc50303a0;  // 0x80000a90
        rom_data[ 677] = 32'h7de20044;  // 0x80000a94
        rom_data[ 678] = 32'hbbe52989;  // 0x80000a98
        rom_data[ 679] = 32'h03000793;  // 0x80000a9c
        rom_data[ 680] = 32'h00f11823;  // 0x80000aa0
        rom_data[ 681] = 32'h08004d05;  // 0x80000aa4
        rom_data[ 682] = 32'h0793b7d1;  // 0x80000aa8
        rom_data[ 683] = 32'h053b02d0;  // 0x80000aac
        rom_data[ 684] = 32'h462940a0;  // 0x80000ab0
        rom_data[ 685] = 32'h01110593;  // 0x80000ab4
        rom_data[ 686] = 32'h00f10823;  // 0x80000ab8
        rom_data[ 687] = 32'hccdff0ef;  // 0x80000abc
        rom_data[ 688] = 32'h00150d1b;  // 0x80000ac0
        rom_data[ 689] = 32'hb75d0800;  // 0x80000ac4
        rom_data[ 690] = 32'h10100713;  // 0x80000ac8
        rom_data[ 691] = 32'h77931742;  // 0x80000acc
        rom_data[ 692] = 32'h8fd90ff5;  // 0x80000ad0
        rom_data[ 693] = 32'h00002717;  // 0x80000ad4
        rom_data[ 694] = 32'h72c70713;  // 0x80000ad8
        rom_data[ 695] = 32'h631ce31c;  // 0x80000adc
        rom_data[ 696] = 32'h8082fffd;  // 0x80000ae0
        rom_data[ 697] = 32'h00054783;  // 0x80000ae4
        rom_data[ 698] = 32'h0613cf8d;  // 0x80000ae8
        rom_data[ 699] = 32'h16421010;  // 0x80000aec
        rom_data[ 700] = 32'h27174681;  // 0x80000af0
        rom_data[ 701] = 32'h07130000;  // 0x80000af4
        rom_data[ 702] = 32'h8fd170e7;  // 0x80000af8
        rom_data[ 703] = 32'h631ce31c;  // 0x80000afc
        rom_data[ 704] = 32'h4783fffd;  // 0x80000b00
        rom_data[ 705] = 32'h05050015;  // 0x80000b04
        rom_data[ 706] = 32'h2685c399;  // 0x80000b08
        rom_data[ 707] = 32'h851bb7fd;  // 0x80000b0c
        rom_data[ 708] = 32'h07930026;  // 0x80000b10
        rom_data[ 709] = 32'h17c21010;  // 0x80000b14
        rom_data[ 710] = 32'he31c07a9;  // 0x80000b18
        rom_data[ 711] = 32'hfffd631c;  // 0x80000b1c
        rom_data[ 712] = 32'h45058082;  // 0x80000b20
        rom_data[ 713] = 32'h00002717;  // 0x80000b24
        rom_data[ 714] = 32'h6dc70713;  // 0x80000b28
        rom_data[ 715] = 32'h0000b7dd;  // 0x80000b2c
        rom_data[ 716] = 32'h0a3a7325;  // 0x80000b30
        rom_data[ 717] = 32'h00000000;  // 0x80000b34
        rom_data[ 718] = 32'h00000000;  // 0x80000b38
        rom_data[ 719] = 32'h00000000;  // 0x80000b3c
        rom_data[ 720] = 32'h005b2020;  // 0x80000b40
        rom_data[ 721] = 32'h00000000;  // 0x80000b44
        rom_data[ 722] = 32'h00643325;  // 0x80000b48
        rom_data[ 723] = 32'h00000000;  // 0x80000b4c
        rom_data[ 724] = 32'h0000005d;  // 0x80000b50
        rom_data[ 725] = 32'h00000000;  // 0x80000b54
        rom_data[ 726] = 32'h0000202c;  // 0x80000b58
        rom_data[ 727] = 32'h00000000;  // 0x80000b5c
        rom_data[ 728] = 32'h00753625;  // 0x80000b60
        rom_data[ 729] = 32'h00000000;  // 0x80000b64
        rom_data[ 730] = 32'h00736559;  // 0x80000b68
        rom_data[ 731] = 32'h00000000;  // 0x80000b6c
        rom_data[ 732] = 32'h00006f4e;  // 0x80000b70
        rom_data[ 733] = 32'h00000000;  // 0x80000b74
        rom_data[ 734] = 32'h203d3d3d;  // 0x80000b78
        rom_data[ 735] = 32'h7274614d;  // 0x80000b7c
        rom_data[ 736] = 32'h41207869;  // 0x80000b80
        rom_data[ 737] = 32'h6c656363;  // 0x80000b84
        rom_data[ 738] = 32'h74617265;  // 0x80000b88
        rom_data[ 739] = 32'h5420726f;  // 0x80000b8c
        rom_data[ 740] = 32'h20747365;  // 0x80000b90
        rom_data[ 741] = 32'h74697553;  // 0x80000b94
        rom_data[ 742] = 32'h3d3d2065;  // 0x80000b98
        rom_data[ 743] = 32'h00000a3d;  // 0x80000b9c
        rom_data[ 744] = 32'h74696e49;  // 0x80000ba0
        rom_data[ 745] = 32'h696c6169;  // 0x80000ba4
        rom_data[ 746] = 32'h676e697a;  // 0x80000ba8
        rom_data[ 747] = 32'h74616d20;  // 0x80000bac
        rom_data[ 748] = 32'h20786972;  // 0x80000bb0
        rom_data[ 749] = 32'h65636361;  // 0x80000bb4
        rom_data[ 750] = 32'h6172656c;  // 0x80000bb8
        rom_data[ 751] = 32'h2e726f74;  // 0x80000bbc
        rom_data[ 752] = 32'h00002e2e;  // 0x80000bc0
        rom_data[ 753] = 32'h00000000;  // 0x80000bc4
        rom_data[ 754] = 32'h4f525245;  // 0x80000bc8
        rom_data[ 755] = 32'h46203a52;  // 0x80000bcc
        rom_data[ 756] = 32'h656c6961;  // 0x80000bd0
        rom_data[ 757] = 32'h6f742064;  // 0x80000bd4
        rom_data[ 758] = 32'h696e6920;  // 0x80000bd8
        rom_data[ 759] = 32'h6c616974;  // 0x80000bdc
        rom_data[ 760] = 32'h20657a69;  // 0x80000be0
        rom_data[ 761] = 32'h65636361;  // 0x80000be4
        rom_data[ 762] = 32'h6172656c;  // 0x80000be8
        rom_data[ 763] = 32'h3a726f74;  // 0x80000bec
        rom_data[ 764] = 32'h0a732520;  // 0x80000bf0
        rom_data[ 765] = 32'h00000000;  // 0x80000bf4
        rom_data[ 766] = 32'h65636341;  // 0x80000bf8
        rom_data[ 767] = 32'h6172656c;  // 0x80000bfc
        rom_data[ 768] = 32'h20726f74;  // 0x80000c00
        rom_data[ 769] = 32'h74696e69;  // 0x80000c04
        rom_data[ 770] = 32'h696c6169;  // 0x80000c08
        rom_data[ 771] = 32'h2064657a;  // 0x80000c0c
        rom_data[ 772] = 32'h63637573;  // 0x80000c10
        rom_data[ 773] = 32'h66737365;  // 0x80000c14
        rom_data[ 774] = 32'h796c6c75;  // 0x80000c18
        rom_data[ 775] = 32'h00000a21;  // 0x80000c1c
        rom_data[ 776] = 32'h74696e49;  // 0x80000c20
        rom_data[ 777] = 32'h206c6169;  // 0x80000c24
        rom_data[ 778] = 32'h74617473;  // 0x80000c28
        rom_data[ 779] = 32'h2d207375;  // 0x80000c2c
        rom_data[ 780] = 32'h73754220;  // 0x80000c30
        rom_data[ 781] = 32'h25203a79;  // 0x80000c34
        rom_data[ 782] = 32'h44202c73;  // 0x80000c38
        rom_data[ 783] = 32'h3a656e6f;  // 0x80000c3c
        rom_data[ 784] = 32'h0a732520;  // 0x80000c40
        rom_data[ 785] = 32'h0000000a;  // 0x80000c44
        rom_data[ 786] = 32'h202d2d2d;  // 0x80000c48
        rom_data[ 787] = 32'h6e6e7552;  // 0x80000c4c
        rom_data[ 788] = 32'h20676e69;  // 0x80000c50
        rom_data[ 789] = 32'h74736554;  // 0x80000c54
        rom_data[ 790] = 32'h73614320;  // 0x80000c58
        rom_data[ 791] = 32'h64252065;  // 0x80000c5c
        rom_data[ 792] = 32'h7325203a;  // 0x80000c60
        rom_data[ 793] = 32'h2d2d2d20;  // 0x80000c64
        rom_data[ 794] = 32'h0000000a;  // 0x80000c68
        rom_data[ 795] = 32'h00000000;  // 0x80000c6c
        rom_data[ 796] = 32'h4f525245;  // 0x80000c70
        rom_data[ 797] = 32'h4d203a52;  // 0x80000c74
        rom_data[ 798] = 32'h69727461;  // 0x80000c78
        rom_data[ 799] = 32'h756d2078;  // 0x80000c7c
        rom_data[ 800] = 32'h7069746c;  // 0x80000c80
        rom_data[ 801] = 32'h6163696c;  // 0x80000c84
        rom_data[ 802] = 32'h6e6f6974;  // 0x80000c88
        rom_data[ 803] = 32'h69616620;  // 0x80000c8c
        rom_data[ 804] = 32'h3a64656c;  // 0x80000c90
        rom_data[ 805] = 32'h0a732520;  // 0x80000c94
        rom_data[ 806] = 32'h00000000;  // 0x80000c98
        rom_data[ 807] = 32'h00000000;  // 0x80000c9c
        rom_data[ 808] = 32'h203d3d3d;  // 0x80000ca0
        rom_data[ 809] = 32'h74736554;  // 0x80000ca4
        rom_data[ 810] = 32'h6d755320;  // 0x80000ca8
        rom_data[ 811] = 32'h7972616d;  // 0x80000cac
        rom_data[ 812] = 32'h3d3d3d20;  // 0x80000cb0
        rom_data[ 813] = 32'h00000000;  // 0x80000cb4
        rom_data[ 814] = 32'h61746f54;  // 0x80000cb8
        rom_data[ 815] = 32'h6574206c;  // 0x80000cbc
        rom_data[ 816] = 32'h3a737473;  // 0x80000cc0
        rom_data[ 817] = 32'h0a642520;  // 0x80000cc4
        rom_data[ 818] = 32'h00000000;  // 0x80000cc8
        rom_data[ 819] = 32'h00000000;  // 0x80000ccc
        rom_data[ 820] = 32'h73736150;  // 0x80000cd0
        rom_data[ 821] = 32'h203a6465;  // 0x80000cd4
        rom_data[ 822] = 32'h000a6425;  // 0x80000cd8
        rom_data[ 823] = 32'h00000000;  // 0x80000cdc
        rom_data[ 824] = 32'h6c696146;  // 0x80000ce0
        rom_data[ 825] = 32'h203a6465;  // 0x80000ce4
        rom_data[ 826] = 32'h000a6425;  // 0x80000ce8
        rom_data[ 827] = 32'h00000000;  // 0x80000cec
        rom_data[ 828] = 32'h63637553;  // 0x80000cf0
        rom_data[ 829] = 32'h20737365;  // 0x80000cf4
        rom_data[ 830] = 32'h65746172;  // 0x80000cf8
        rom_data[ 831] = 32'h2e25203a;  // 0x80000cfc
        rom_data[ 832] = 32'h25256631;  // 0x80000d00
        rom_data[ 833] = 32'h0000000a;  // 0x80000d04
        rom_data[ 834] = 32'h8e9ff00a;  // 0x80000d08
        rom_data[ 835] = 32'h6c412089;  // 0x80000d0c
        rom_data[ 836] = 32'h6574206c;  // 0x80000d10
        rom_data[ 837] = 32'h20737473;  // 0x80000d14
        rom_data[ 838] = 32'h73736170;  // 0x80000d18
        rom_data[ 839] = 32'h20216465;  // 0x80000d1c
        rom_data[ 840] = 32'h7274614d;  // 0x80000d20
        rom_data[ 841] = 32'h61207869;  // 0x80000d24
        rom_data[ 842] = 32'h6c656363;  // 0x80000d28
        rom_data[ 843] = 32'h74617265;  // 0x80000d2c
        rom_data[ 844] = 32'h6920726f;  // 0x80000d30
        rom_data[ 845] = 32'h6f772073;  // 0x80000d34
        rom_data[ 846] = 32'h6e696b72;  // 0x80000d38
        rom_data[ 847] = 32'h6f632067;  // 0x80000d3c
        rom_data[ 848] = 32'h63657272;  // 0x80000d40
        rom_data[ 849] = 32'h2e796c74;  // 0x80000d44
        rom_data[ 850] = 32'h00000000;  // 0x80000d48
        rom_data[ 851] = 32'h00000000;  // 0x80000d4c
        rom_data[ 852] = 32'h2d2d2d0a;  // 0x80000d50
        rom_data[ 853] = 32'h6e755220;  // 0x80000d54
        rom_data[ 854] = 32'h676e696e;  // 0x80000d58
        rom_data[ 855] = 32'h72655020;  // 0x80000d5c
        rom_data[ 856] = 32'h6d726f66;  // 0x80000d60
        rom_data[ 857] = 32'h65636e61;  // 0x80000d64
        rom_data[ 858] = 32'h73655420;  // 0x80000d68
        rom_data[ 859] = 32'h2d2d2074;  // 0x80000d6c
        rom_data[ 860] = 32'h0000002d;  // 0x80000d70
        rom_data[ 861] = 32'h00000000;  // 0x80000d74
        rom_data[ 862] = 32'h6e6e7552;  // 0x80000d78
        rom_data[ 863] = 32'h20676e69;  // 0x80000d7c
        rom_data[ 864] = 32'h66726570;  // 0x80000d80
        rom_data[ 865] = 32'h616d726f;  // 0x80000d84
        rom_data[ 866] = 32'h2065636e;  // 0x80000d88
        rom_data[ 867] = 32'h74736574;  // 0x80000d8c
        rom_data[ 868] = 32'h74697720;  // 0x80000d90
        rom_data[ 869] = 32'h616c2068;  // 0x80000d94
        rom_data[ 870] = 32'h72656772;  // 0x80000d98
        rom_data[ 871] = 32'h6c617620;  // 0x80000d9c
        rom_data[ 872] = 32'h2e736575;  // 0x80000da0
        rom_data[ 873] = 32'h00002e2e;  // 0x80000da4
        rom_data[ 874] = 32'h66726550;  // 0x80000da8
        rom_data[ 875] = 32'h616d726f;  // 0x80000dac
        rom_data[ 876] = 32'h2065636e;  // 0x80000db0
        rom_data[ 877] = 32'h7274614d;  // 0x80000db4
        rom_data[ 878] = 32'h41207869;  // 0x80000db8
        rom_data[ 879] = 32'h00000000;  // 0x80000dbc
        rom_data[ 880] = 32'h66726550;  // 0x80000dc0
        rom_data[ 881] = 32'h616d726f;  // 0x80000dc4
        rom_data[ 882] = 32'h2065636e;  // 0x80000dc8
        rom_data[ 883] = 32'h7274614d;  // 0x80000dcc
        rom_data[ 884] = 32'h42207869;  // 0x80000dd0
        rom_data[ 885] = 32'h00000000;  // 0x80000dd4
        rom_data[ 886] = 32'h66726550;  // 0x80000dd8
        rom_data[ 887] = 32'h616d726f;  // 0x80000ddc
        rom_data[ 888] = 32'h2065636e;  // 0x80000de0
        rom_data[ 889] = 32'h74736574;  // 0x80000de4
        rom_data[ 890] = 32'h6d6f6320;  // 0x80000de8
        rom_data[ 891] = 32'h74656c70;  // 0x80000dec
        rom_data[ 892] = 32'h73206465;  // 0x80000df0
        rom_data[ 893] = 32'h65636375;  // 0x80000df4
        rom_data[ 894] = 32'h75667373;  // 0x80000df8
        rom_data[ 895] = 32'h21796c6c;  // 0x80000dfc
        rom_data[ 896] = 32'h00000000;  // 0x80000e00
        rom_data[ 897] = 32'h00000000;  // 0x80000e04
        rom_data[ 898] = 32'h66726550;  // 0x80000e08
        rom_data[ 899] = 32'h616d726f;  // 0x80000e0c
        rom_data[ 900] = 32'h2065636e;  // 0x80000e10
        rom_data[ 901] = 32'h75736552;  // 0x80000e14
        rom_data[ 902] = 32'h0000746c;  // 0x80000e18
        rom_data[ 903] = 32'h00000000;  // 0x80000e1c
        rom_data[ 904] = 32'h69747345;  // 0x80000e20
        rom_data[ 905] = 32'h6574616d;  // 0x80000e24
        rom_data[ 906] = 32'h79632064;  // 0x80000e28
        rom_data[ 907] = 32'h73656c63;  // 0x80000e2c
        rom_data[ 908] = 32'h7525203a;  // 0x80000e30
        rom_data[ 909] = 32'h0000000a;  // 0x80000e34
        rom_data[ 910] = 32'h65746f4e;  // 0x80000e38
        rom_data[ 911] = 32'h7943203a;  // 0x80000e3c
        rom_data[ 912] = 32'h20656c63;  // 0x80000e40
        rom_data[ 913] = 32'h6e756f63;  // 0x80000e44
        rom_data[ 914] = 32'h676e6974;  // 0x80000e48
        rom_data[ 915] = 32'h746f6e20;  // 0x80000e4c
        rom_data[ 916] = 32'h706d6920;  // 0x80000e50
        rom_data[ 917] = 32'h656d656c;  // 0x80000e54
        rom_data[ 918] = 32'h6465746e;  // 0x80000e58
        rom_data[ 919] = 32'h206e6920;  // 0x80000e5c
        rom_data[ 920] = 32'h73696874;  // 0x80000e60
        rom_data[ 921] = 32'h73657420;  // 0x80000e64
        rom_data[ 922] = 32'h65762074;  // 0x80000e68
        rom_data[ 923] = 32'h6f697372;  // 0x80000e6c
        rom_data[ 924] = 32'h0000006e;  // 0x80000e70
        rom_data[ 925] = 32'h00000000;  // 0x80000e74
        rom_data[ 926] = 32'h66726550;  // 0x80000e78
        rom_data[ 927] = 32'h616d726f;  // 0x80000e7c
        rom_data[ 928] = 32'h2065636e;  // 0x80000e80
        rom_data[ 929] = 32'h74736574;  // 0x80000e84
        rom_data[ 930] = 32'h69616620;  // 0x80000e88
        rom_data[ 931] = 32'h3a64656c;  // 0x80000e8c
        rom_data[ 932] = 32'h0a732520;  // 0x80000e90
        rom_data[ 933] = 32'h00000000;  // 0x80000e94
        rom_data[ 934] = 32'h8c9de20a;  // 0x80000e98
        rom_data[ 935] = 32'h6d6f5320;  // 0x80000e9c
        rom_data[ 936] = 32'h65742065;  // 0x80000ea0
        rom_data[ 937] = 32'h20737473;  // 0x80000ea4
        rom_data[ 938] = 32'h6c696166;  // 0x80000ea8
        rom_data[ 939] = 32'h202e6465;  // 0x80000eac
        rom_data[ 940] = 32'h61656c50;  // 0x80000eb0
        rom_data[ 941] = 32'h63206573;  // 0x80000eb4
        rom_data[ 942] = 32'h6b636568;  // 0x80000eb8
        rom_data[ 943] = 32'h65687420;  // 0x80000ebc
        rom_data[ 944] = 32'h72616820;  // 0x80000ec0
        rom_data[ 945] = 32'h72617764;  // 0x80000ec4
        rom_data[ 946] = 32'h6d692065;  // 0x80000ec8
        rom_data[ 947] = 32'h6d656c70;  // 0x80000ecc
        rom_data[ 948] = 32'h61746e65;  // 0x80000ed0
        rom_data[ 949] = 32'h6e6f6974;  // 0x80000ed4
        rom_data[ 950] = 32'h0000002e;  // 0x80000ed8
        rom_data[ 951] = 32'h00000000;  // 0x80000edc
        rom_data[ 952] = 32'h53534150;  // 0x80000ee0
        rom_data[ 953] = 32'h6554203a;  // 0x80000ee4
        rom_data[ 954] = 32'h63207473;  // 0x80000ee8
        rom_data[ 955] = 32'h20657361;  // 0x80000eec
        rom_data[ 956] = 32'h70206425;  // 0x80000ef0
        rom_data[ 957] = 32'h65737361;  // 0x80000ef4
        rom_data[ 958] = 32'h000a2164;  // 0x80000ef8
        rom_data[ 959] = 32'h00000000;  // 0x80000efc
        rom_data[ 960] = 32'h4c494146;  // 0x80000f00
        rom_data[ 961] = 32'h6554203a;  // 0x80000f04
        rom_data[ 962] = 32'h63207473;  // 0x80000f08
        rom_data[ 963] = 32'h20657361;  // 0x80000f0c
        rom_data[ 964] = 32'h66206425;  // 0x80000f10
        rom_data[ 965] = 32'h656c6961;  // 0x80000f14
        rom_data[ 966] = 32'h000a2164;  // 0x80000f18
        rom_data[ 967] = 32'h00000000;  // 0x80000f1c
        rom_data[ 968] = 32'h7274614d;  // 0x80000f20
        rom_data[ 969] = 32'h41207869;  // 0x80000f24
        rom_data[ 970] = 32'h00000000;  // 0x80000f28
        rom_data[ 971] = 32'h00000000;  // 0x80000f2c
        rom_data[ 972] = 32'h7274614d;  // 0x80000f30
        rom_data[ 973] = 32'h42207869;  // 0x80000f34
        rom_data[ 974] = 32'h00000000;  // 0x80000f38
        rom_data[ 975] = 32'h00000000;  // 0x80000f3c
        rom_data[ 976] = 32'h65707845;  // 0x80000f40
        rom_data[ 977] = 32'h64657463;  // 0x80000f44
        rom_data[ 978] = 32'h00000000;  // 0x80000f48
        rom_data[ 979] = 32'h00000000;  // 0x80000f4c
        rom_data[ 980] = 32'h75746341;  // 0x80000f50
        rom_data[ 981] = 32'h00006c61;  // 0x80000f54
        rom_data[ 982] = 32'h6e656449;  // 0x80000f58
        rom_data[ 983] = 32'h79746974;  // 0x80000f5c
        rom_data[ 984] = 32'h74614d20;  // 0x80000f60
        rom_data[ 985] = 32'h20786972;  // 0x80000f64
        rom_data[ 986] = 32'h74736554;  // 0x80000f68
        rom_data[ 987] = 32'h00000000;  // 0x80000f6c
        rom_data[ 988] = 32'h706d6953;  // 0x80000f70
        rom_data[ 989] = 32'h4d20656c;  // 0x80000f74
        rom_data[ 990] = 32'h69746c75;  // 0x80000f78
        rom_data[ 991] = 32'h63696c70;  // 0x80000f7c
        rom_data[ 992] = 32'h6f697461;  // 0x80000f80
        rom_data[ 993] = 32'h6554206e;  // 0x80000f84
        rom_data[ 994] = 32'h00007473;  // 0x80000f88
        rom_data[ 995] = 32'h00000000;  // 0x80000f8c
        rom_data[ 996] = 32'h206c6c41;  // 0x80000f90
        rom_data[ 997] = 32'h73656e4f;  // 0x80000f94
        rom_data[ 998] = 32'h73655420;  // 0x80000f98
        rom_data[ 999] = 32'h00000074;  // 0x80000f9c
        rom_data[1000] = 32'h6e6b6e55;  // 0x80000fa0
        rom_data[1001] = 32'h206e776f;  // 0x80000fa4
        rom_data[1002] = 32'h6f727265;  // 0x80000fa8
        rom_data[1003] = 32'h00000072;  // 0x80000fac
        rom_data[1004] = 32'h61766e49;  // 0x80000fb0
        rom_data[1005] = 32'h2064696c;  // 0x80000fb4
        rom_data[1006] = 32'h61726170;  // 0x80000fb8
        rom_data[1007] = 32'h6574656d;  // 0x80000fbc
        rom_data[1008] = 32'h00000072;  // 0x80000fc0
        rom_data[1009] = 32'h00000000;  // 0x80000fc4
        rom_data[1010] = 32'h65636341;  // 0x80000fc8
        rom_data[1011] = 32'h6172656c;  // 0x80000fcc
        rom_data[1012] = 32'h20726f74;  // 0x80000fd0
        rom_data[1013] = 32'h79737562;  // 0x80000fd4
        rom_data[1014] = 32'h00000000;  // 0x80000fd8
        rom_data[1015] = 32'h00000000;  // 0x80000fdc
        rom_data[1016] = 32'h7265704f;  // 0x80000fe0
        rom_data[1017] = 32'h6f697461;  // 0x80000fe4
        rom_data[1018] = 32'h6974206e;  // 0x80000fe8
        rom_data[1019] = 32'h756f656d;  // 0x80000fec
        rom_data[1020] = 32'h00000074;  // 0x80000ff0
        rom_data[1021] = 32'h00000000;  // 0x80000ff4
        rom_data[1022] = 32'h63637553;  // 0x80000ff8
        rom_data[1023] = 32'h00737365;  // 0x80000ffc
        rom_data[1024] = 32'h33323130;  // 0x80001000
        rom_data[1025] = 32'h37363534;  // 0x80001004
        rom_data[1026] = 32'h42413938;  // 0x80001008
        rom_data[1027] = 32'h46454443;  // 0x8000100c
        rom_data[1028] = 32'h00000000;  // 0x80001010
        rom_data[1029] = 32'h00000000;  // 0x80001014
        rom_data[1030] = 32'h80000f58;  // 0x80001018
        rom_data[1031] = 32'h00000000;  // 0x8000101c
        rom_data[1032] = 32'h04030201;  // 0x80001020
        rom_data[1033] = 32'h08070605;  // 0x80001024
        rom_data[1034] = 32'h0c0b0a09;  // 0x80001028
        rom_data[1035] = 32'h100f0e0d;  // 0x8000102c
        rom_data[1036] = 32'h00000001;  // 0x80001030
        rom_data[1037] = 32'h00000100;  // 0x80001034
        rom_data[1038] = 32'h00010000;  // 0x80001038
        rom_data[1039] = 32'h01000000;  // 0x8000103c
        rom_data[1040] = 32'h00000001;  // 0x80001040
        rom_data[1041] = 32'h00000002;  // 0x80001044
        rom_data[1042] = 32'h00000003;  // 0x80001048
        rom_data[1043] = 32'h00000004;  // 0x8000104c
        rom_data[1044] = 32'h00000005;  // 0x80001050
        rom_data[1045] = 32'h00000006;  // 0x80001054
        rom_data[1046] = 32'h00000007;  // 0x80001058
        rom_data[1047] = 32'h00000008;  // 0x8000105c
        rom_data[1048] = 32'h00000009;  // 0x80001060
        rom_data[1049] = 32'h0000000a;  // 0x80001064
        rom_data[1050] = 32'h0000000b;  // 0x80001068
        rom_data[1051] = 32'h0000000c;  // 0x8000106c
        rom_data[1052] = 32'h0000000d;  // 0x80001070
        rom_data[1053] = 32'h0000000e;  // 0x80001074
        rom_data[1054] = 32'h0000000f;  // 0x80001078
        rom_data[1055] = 32'h00000010;  // 0x8000107c
        rom_data[1056] = 32'h80000f70;  // 0x80001080
        rom_data[1057] = 32'h00000000;  // 0x80001084
        rom_data[1058] = 32'h00000201;  // 0x80001088
        rom_data[1059] = 32'h00020100;  // 0x8000108c
        rom_data[1060] = 32'h02010000;  // 0x80001090
        rom_data[1061] = 32'h01000000;  // 0x80001094
        rom_data[1062] = 32'h00000002;  // 0x80001098
        rom_data[1063] = 32'h00000201;  // 0x8000109c
        rom_data[1064] = 32'h00020100;  // 0x800010a0
        rom_data[1065] = 32'h02010000;  // 0x800010a4
        rom_data[1066] = 32'h00000004;  // 0x800010a8
        rom_data[1067] = 32'h00000004;  // 0x800010ac
        rom_data[1068] = 32'h00000000;  // 0x800010b0
        rom_data[1069] = 32'h00000000;  // 0x800010b4
        rom_data[1070] = 32'h00000001;  // 0x800010b8
        rom_data[1071] = 32'h00000004;  // 0x800010bc
        rom_data[1072] = 32'h00000004;  // 0x800010c0
        rom_data[1073] = 32'h00000000;  // 0x800010c4
        rom_data[1074] = 32'h00000000;  // 0x800010c8
        rom_data[1075] = 32'h00000001;  // 0x800010cc
        rom_data[1076] = 32'h00000004;  // 0x800010d0
        rom_data[1077] = 32'h00000004;  // 0x800010d4
        rom_data[1078] = 32'h00000000;  // 0x800010d8
        rom_data[1079] = 32'h00000000;  // 0x800010dc
        rom_data[1080] = 32'h00000001;  // 0x800010e0
        rom_data[1081] = 32'h00000002;  // 0x800010e4
        rom_data[1082] = 32'h80000f90;  // 0x800010e8
        rom_data[1083] = 32'h00000000;  // 0x800010ec
        rom_data[1084] = 32'h01010101;  // 0x800010f0
        rom_data[1085] = 32'h01010101;  // 0x800010f4
        rom_data[1086] = 32'h01010101;  // 0x800010f8
        rom_data[1087] = 32'h01010101;  // 0x800010fc
        rom_data[1088] = 32'h01010101;  // 0x80001100
        rom_data[1089] = 32'h01010101;  // 0x80001104
        rom_data[1090] = 32'h01010101;  // 0x80001108
        rom_data[1091] = 32'h01010101;  // 0x8000110c
        rom_data[1092] = 32'h00000004;  // 0x80001110
        rom_data[1093] = 32'h00000004;  // 0x80001114
        rom_data[1094] = 32'h00000004;  // 0x80001118
        rom_data[1095] = 32'h00000004;  // 0x8000111c
        rom_data[1096] = 32'h00000004;  // 0x80001120
        rom_data[1097] = 32'h00000004;  // 0x80001124
        rom_data[1098] = 32'h00000004;  // 0x80001128
        rom_data[1099] = 32'h00000004;  // 0x8000112c
        rom_data[1100] = 32'h00000004;  // 0x80001130
        rom_data[1101] = 32'h00000004;  // 0x80001134
        rom_data[1102] = 32'h00000004;  // 0x80001138
        rom_data[1103] = 32'h00000004;  // 0x8000113c
        rom_data[1104] = 32'h00000004;  // 0x80001140
        rom_data[1105] = 32'h00000004;  // 0x80001144
        rom_data[1106] = 32'h00000004;  // 0x80001148
        rom_data[1107] = 32'h00000004;  // 0x8000114c
        rom_data[1108] = 32'h281e140a;  // 0x80001150
        rom_data[1109] = 32'h50463c32;  // 0x80001154
        rom_data[1110] = 32'h786e645a;  // 0x80001158
        rom_data[1111] = 32'ha0968c82;  // 0x8000115c
        rom_data[1112] = 32'h04030201;  // 0x80001160
        rom_data[1113] = 32'h08070605;  // 0x80001164
        rom_data[1114] = 32'h0c0b0a09;  // 0x80001168
        rom_data[1115] = 32'h100f0e0d;  // 0x8000116c
        rom_data[1116] = 32'h80000fb0;  // 0x80001170
        rom_data[1117] = 32'h00000000;  // 0x80001174
        rom_data[1118] = 32'h80000fc8;  // 0x80001178
        rom_data[1119] = 32'h00000000;  // 0x8000117c
        rom_data[1120] = 32'h80000fe0;  // 0x80001180
        rom_data[1121] = 32'h00000000;  // 0x80001184
        rom_data[1122] = 32'h80000ff8;  // 0x80001188
        rom_data[1123] = 32'h00000000;  // 0x8000118c
        rom_data[1124] = 32'hfffff7f6;  // 0x80001190
        rom_data[1125] = 32'hfffff7be;  // 0x80001194
        rom_data[1126] = 32'hfffff6ec;  // 0x80001198
        rom_data[1127] = 32'hfffff6ec;  // 0x8000119c
        rom_data[1128] = 32'hfffff6ec;  // 0x800011a0
        rom_data[1129] = 32'hfffff6ec;  // 0x800011a4
        rom_data[1130] = 32'hfffff6ec;  // 0x800011a8
        rom_data[1131] = 32'hfffff6ec;  // 0x800011ac
        rom_data[1132] = 32'hfffff6ec;  // 0x800011b0
        rom_data[1133] = 32'hfffff6ec;  // 0x800011b4
        rom_data[1134] = 32'hfffff6ec;  // 0x800011b8
        rom_data[1135] = 32'hfffff6ec;  // 0x800011bc
        rom_data[1136] = 32'hfffff6ec;  // 0x800011c0
        rom_data[1137] = 32'hfffff6ec;  // 0x800011c4
        rom_data[1138] = 32'hfffff6ec;  // 0x800011c8
        rom_data[1139] = 32'hfffff6ec;  // 0x800011cc
        rom_data[1140] = 32'hfffff792;  // 0x800011d0
        rom_data[1141] = 32'hfffff6ec;  // 0x800011d4
        rom_data[1142] = 32'hfffff75c;  // 0x800011d8
        rom_data[1143] = 32'hfffff6ec;  // 0x800011dc
        rom_data[1144] = 32'hfffff6ec;  // 0x800011e0
        rom_data[1145] = 32'hfffff726;  // 0x800011e4
        rom_data[1146] = 32'h40400000;  // 0x800011e8
        rom_data[1147] = 32'h42c80000;  // 0x800011ec
        rom_data[1148] = 32'h00000000;  // 0x800011f0
        rom_data[1149] = 32'h40240000;  // 0x800011f4
    end

endmodule
